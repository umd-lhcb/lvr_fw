--------------------------------------------------------------------------------
-- Company: UNIVERSITY OF MARYLAND
--
-- File: SERIAL_TX.vhd
-- File history:
--      <Rev - // Mar 30, 2017  INITIAL
--
-- Description: THIS MODULE TRANSMITS THE SERIAL WORD.
--					FRAME PACKET CONSISTS OF 16 BITS + 2 START AND 2 STOP BITS.
--					LSB ASSUMED FIRST
--					THE START AND STOP BITS ARE ALL LOGIC '1'----!!!! THE STOP BIT NEEDS TO BE FOLLOWED BY A FORCED '0' !!!!!!
--					15		ODD PARITY (APPLIES TO 15 DATA BITS ONLY (14:0) )
--					14		UVL STATUS
--					13..12	MODE 
--					11..8	MODULE ADDRESS
--					7..0	CHANNEL ENABLES
--					
--					
--					BIT IS DERIVED FROM 5 MHZ CLOCK DIVIDED BY 64 = 12.8 USEC (78.125 KBPS)
--					12.8 USEC / 200NS = 64 COUNTS
--
--
-- Targeted device: <Family::ProASIC3> <Die::A3PN125> <Package::100 VQFP>
-- Author: TOM O'BANNON
--
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_MISC.ALL;
USE IEEE.NUMERIC_STD.ALL;

library proasic3;
use proasic3.all;

-- NOTE:  THE SYNPLIFY LIBRARY NEEDS TO BE COMMENTED OUT FOR MODELSIM PRESYNTH SIMS SINCE MODELSIM DOES NOT RECOGNIZE IT
library synplify;
use synplify.attributes.all;

entity SERIAL_TX is
port (
		MASTER_RST_B		:	IN	STD_LOGIC;							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
		CLK_5M_GL			:	IN	STD_LOGIC;
		TX_WORD				:	IN	STD_LOGIC_VECTOR(14 DOWNTO 0);		-- PARALLEL WORD TO BE TRANSMITTED (NOTE--BIT 15 IS ODD PARITY CALCULATED AS SERIAL TX IS SENT)
		TX_STRB				:	IN	STD_LOGIC;							-- SINGLE CLOCK PULSE STRB INDICATES NEW TX_WORD READY FOR TX
		
		P_TX_EN				:	OUT	STD_LOGIC;							-- SERIAL TX DRIVER ENABLE
		SER_TX_BIT			:	OUT	STD_LOGIC							-- TX BIT STREAM
	);
end SERIAL_TX;

architecture RTL of SERIAL_TX is
ATTRIBUTE SYN_RADHARDLEVEL OF RTL : ARCHITECTURE IS "TMR";

-- !!!!!  NOTE   !!!! THE STATE MACHINES NEED TO HAVE THE "SAFE ATTRIBUTE" APPLIED IN SYNTHESIS

-- DEFINE THE STATES FOR SERIAL RECEIVE STATE MACHINE-----!!!!! ADD PLACEHOLDERS TO CREATE 2^^N STATES !!!!!!
TYPE TRANSMIT_STATES IS (	INIT, BIT_DEL_WAIT, TX_1ST_START_BIT, TX_2ND_START_BIT, 
					TX_0LS_BIT, TX_1_BIT, TX_2_BIT, TX_3_BIT, TX_4_BIT, TX_5_BIT, TX_6_BIT, TX_7_BIT, 
					TX_8_BIT, TX_9_BIT, TX_10_BIT, TX_11_BIT, TX_12_BIT, TX_13_BIT, TX_14_BIT, TX_15_BIT, 
					TX_1ST_STOP_BIT, TX_2ND_STOP_BIT, FINISH_FRAME, FINISH_STROBE
					);

SIGNAL 	N_TX_STATE, TX_STATE 				: 	TRANSMIT_STATES;							-- STATE MACHINE COUNTER FOR THE RX STATE MACHINE
SIGNAL	N_RET_STATE, RET_STATE				:	TRANSMIT_STATES;							-- POINTER FOR A RETURN LOCATION ON THE RX STATE MACHINE

SIGNAL	N_BIT_POSN_CNT, BIT_POSN_CNT		:	INTEGER RANGE 0 TO 127;						-- COUNTER USED TO MEASURE BIT POSITION EVENTS
SIGNAL	N_TX_BIT, TX_BIT					:	STD_LOGIC;									-- TX SERIAL BIT BUFFER
SIGNAL  N_TX_EN, TX_EN						:	STD_LOGIC;									-- TX DRIVER ENABLE
SIGNAL	N_ODD_PARITY, ODD_PARITY			:	STD_LOGIC;									-- ODD PARITY BIT FOR RX WORD

CONSTANT 	FULL_BIT_CNT					:	INTEGER RANGE 0 TO 127 := 61;				-- 64 COUNTS OF 5 MHZ CLOCK = FULL SERIAL BIT POSITION, 
																							-- BUT NEED 2 LESS TO ALLOW FOR STATE MACHINE STEPS IN AND OUT OF BIT COUNTER STATE

begin

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE ALL REGISTERS USED WITH THE 5 MHZ CLOCK
REG5M:PROCESS(CLK_5M_GL, MASTER_RST_B)	
	BEGIN
		IF MASTER_RST_B = '0' THEN
			TX_STATE		<=	INIT;
			BIT_POSN_CNT	<=	 0;
			TX_BIT			<=	'0';
			TX_EN			<=	'0';
			ODD_PARITY		<=	'0';
			RET_STATE		<=	INIT;
			
		ELSIF (CLK_5M_GL'EVENT AND CLK_5M_GL='1') THEN
			TX_STATE		<=	N_TX_STATE;
			BIT_POSN_CNT	<=	N_BIT_POSN_CNT;
			TX_BIT			<=	N_TX_BIT;
			TX_EN			<=	N_TX_EN	;
			ODD_PARITY		<=	N_ODD_PARITY;
			RET_STATE		<=	N_RET_STATE;
			
		END IF;
		
	END PROCESS;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE THE SERIAL RX PROCESS
SER_RX:PROCESS(TX_STATE, RET_STATE, BIT_POSN_CNT, TX_WORD, TX_STRB, TX_BIT, TX_EN, ODD_PARITY)
	BEGIN
	
	-- DEFAULT ASSIGNMENTS (GET OVER-WRITTEN BELOW AS NEEDED)
	N_RET_STATE			<=	RET_STATE;
	N_BIT_POSN_CNT		<=	BIT_POSN_CNT;
	N_ODD_PARITY		<=	ODD_PARITY;
	N_TX_BIT			<=	TX_BIT;
	N_TX_EN				<=	TX_EN;
	
		CASE TX_STATE IS

			WHEN INIT			=>									-- WAIT HERE FOR A LOGIC 1 DETECTION ON THE TX_STRB
				IF TX_STRB = '1'	THEN
					N_TX_STATE		<=	TX_1ST_START_BIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
					N_TX_EN			<=	'1';						-- ENABLE THE TRANSMIT SERIAL DRIVER
				ELSE
					N_TX_STATE		<=	INIT;						-- STAY HERE UNLESS '1' DETECTED ON TX_STRB
					N_TX_EN			<=	'0';						-- DISABLE THE TRANSMIT SERIAL DRIVER
				END IF;

				N_ODD_PARITY	<=	 '0';							-- INITIALIZE THE TX ODD PARITY BIT

			WHEN BIT_DEL_WAIT	=>									-- WAIT HERE FOR THE SPECIFIED BIT TIME DELAY--THIS STATE STEP IS REUSED TO MEASURE EACH 1 BIT DURATION
				IF  BIT_POSN_CNT = 0	THEN
					N_TX_STATE		<=	RET_STATE;					-- BRANCH TO THE NEXT STATE
					N_BIT_POSN_CNT	<=	FULL_BIT_CNT;				-- REINITIALIZE FOR THE FULL BIT COUNT VALUE
				ELSE
					N_TX_STATE		<=	BIT_DEL_WAIT;				-- STAY HERE UNTIL DONE
					N_BIT_POSN_CNT	<=	BIT_POSN_CNT - 1;			-- DECREMENT THE COUNTER
				END IF;
				
			WHEN TX_1ST_START_BIT	=>								-- TRANSMIT THE FIRST START BIT
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_2ND_START_BIT;			-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_TX_BIT			<=	'1';
				
			WHEN TX_2ND_START_BIT	=>								-- TRANSMIT THE SECOND START BIT
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_0LS_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_TX_BIT			<=	'1';

			WHEN TX_0LS_BIT			=>								-- TRANSMIT THE LSB 0 BIT VALUE
				N_TX_BIT			<=	TX_WORD(0);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_1_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(0);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_1_BIT		=>									-- TRANSMIT THE BIT 1 VALUE
				N_TX_BIT			<=	TX_WORD(1);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_2_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(1);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_2_BIT		=>									-- TRANSMIT THE BIT 2 VALUE
				N_TX_BIT			<=	TX_WORD(2);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_3_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(2);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_3_BIT		=>									-- TRANSMIT THE BIT 3 VALUE
				N_TX_BIT			<=	TX_WORD(3);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_4_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(3);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_4_BIT		=>									-- TRANSMIT THE BIT 4 VALUE
				N_TX_BIT			<=	TX_WORD(4);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_5_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(4);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_5_BIT		=>									-- TRANSMIT THE BIT 5 VALUE
				N_TX_BIT			<=	TX_WORD(5);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_6_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(5);	-- CALCULATE THE RUNNING PARITY
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE

			WHEN TX_6_BIT		=>									-- TRANSMIT THE BIT 6 VALUE
				N_TX_BIT			<=	TX_WORD(6);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_7_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(6);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_7_BIT		=>									-- TRANSMIT THE BIT 7 VALUE
				N_TX_BIT			<=	TX_WORD(7);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_8_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(7);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_8_BIT		=>									-- TRANSMIT THE BIT 8 VALUE
				N_TX_BIT			<=	TX_WORD(8);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_9_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(8);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_9_BIT		=>									-- TRANSMIT THE BIT 9 VALUE
				N_TX_BIT			<=	TX_WORD(9);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_10_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(9);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_10_BIT		=>									-- TRANSMIT THE BIT 10 VALUE
				N_TX_BIT			<=	TX_WORD(10);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_11_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(10);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_11_BIT		=>									-- TRANSMIT THE BIT 11 VALUE
				N_TX_BIT			<=	TX_WORD(11);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_12_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(11);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_12_BIT		=>									-- TRANSMIT THE BIT 12 VALUE
				N_TX_BIT			<=	TX_WORD(12);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_13_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(12);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_13_BIT		=>									-- TRANSMIT THE BIT 13 VALUE
				N_TX_BIT			<=	TX_WORD(13);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_14_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(13);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_14_BIT		=>									-- TRANSMIT THE BIT 14 VALUE
				N_TX_BIT			<=	TX_WORD(14);
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_15_BIT;					-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR TX_WORD(14);	-- CALCULATE THE RUNNING PARITY

			WHEN TX_15_BIT		=>									-- TRANSMIT THE BIT 15 VALUE WHICH IS THE ODD PARITY FOR THE PREVIOUS 15 DATA BITS
				N_TX_BIT			<=	ODD_PARITY;
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_1ST_STOP_BIT;			-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				
			WHEN TX_1ST_STOP_BIT	=>								-- TRANSMIT THE FIRST STOP BIT
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	TX_2ND_STOP_BIT;			-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_TX_BIT			<=	'1';
				
			WHEN TX_2ND_STOP_BIT	=>								-- TRANSMIT THE SECOND STOP BIT
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	FINISH_FRAME;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_TX_BIT			<=	'1';
			
			WHEN FINISH_FRAME	=>									-- LEAVE THE TX SERIAL OUTPUT IN ZERO POSITION FOR 1 BIT DURATION (THEN MASTER TX NEEDS TO CONTINUE ASSERTING A '0')
				N_TX_STATE			<=	BIT_DEL_WAIT;				-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	FINISH_STROBE;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;				-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_TX_BIT			<=	'0';

			WHEN FINISH_STROBE		=>	
				N_TX_STATE			<=	INIT;						-- 			
				N_TX_BIT			<=	'0';						-- LEAVE THE OUTPUT BIT AT ZERO TO AVOID ANOTHER START BIT DETECTION BY A SERIAL RECEIVER
				N_TX_EN				<=	'0';						-- DISABLE THE TRANSMIT SERIAL DRIVER
			
		END CASE;

	END PROCESS;
	
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- ASSIGN INTERNAL SIGNALS TO EXTERNAL PORTS 
SER_TX_BIT		<=	TX_BIT;
P_TX_EN			<=	TX_EN;
	
end RTL;
