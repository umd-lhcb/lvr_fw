--------------------------------------------------------------------------------
-- Company: University of Maryland
--
-- File: SPI_ALT.vhd
-- File history:
--      INIT, APRIL 3, 2019
--      
--
-- Description: 
--
-- SPI PORT: 	SLAVE IMPLEMENTATION WITHOUT USING SLAVE SELECTS
--				NOTE:  THE CLOCK FOR THE INTERFACE ORIGINATES FROM THE SCA MASTER IN ALL DATA EXCHANGES
--				DATA RATE = 312.5 Kbps (IE ACTUAL SERIAL CLOCK FREQUENCY = LHC 40MHZ / 128 )
--					
-- 	SCA_CLK_OUT		:  	CLOCK INPUT TO THE FPGA FROM THE SCA MASTER
-- 	SCA_DAT_IN		:	DATA OUTPUT FROM THE FPGA TO THE SCA MASTER
-- 	SCA_DAT_OUT		:	DATA INPUT TO THE FPGA FROM THE SCA MASTER
--
-- Targeted device: <Family::ProASIC3> <Die::A3PN250> <Package::100 VQFP>
-- Author: Tom O'Bannon
--
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_MISC.ALL;
--USE IEEE.NUMERIC_STD.ALL;

library proasic3;
use proasic3.all;
	
entity SPI_alt is
port (
        CLK5M_OSC          		:   IN  STD_LOGIC;                      	-- INTERNAL GENERATED 5 MHZ CLOCK 
        MASTER_RST_B           	:   IN  STD_LOGIC;                         	-- INTERNAL ACTIVE LOW RESET

		SCA_CLK_OUT				:  	IN	STD_LOGIC;							-- CLOCK INPUT TO THE FPGA FROM THE SCA MASTER USED FOR BOTH TX AND RX
		SCA_DAT_OUT				:	IN	STD_LOGIC;							-- SERIAL DATA INPUT TO THE FPGA FROM THE SCA MASTER
		SCA_DAT_IN				:	OUT	STD_LOGIC;							-- SERIAL DATA OUTPUT FROM THE FPGA TO THE SCA MASTER

		SPI_TX_WORD				:	IN 	STD_LOGIC_VECTOR(31 DOWNTO 0);		-- 32 BIT SERIAL WORD TO BE TRANSMITTED
		SPI_RX_WORD				:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);		-- RECEIVED SERIAL FRAME
		SPI_RX_STRB				:	OUT	STD_LOGIC;							-- SINGLE 5MHZ CLOCK PULSE SIGNIFIES A NEW SERIAL FRAME IS AVAILABLE.

		P_TX_32BIT_REG			:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		P_STATE_ID				:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0)

	);
end SPI_ALT;

architecture RTL of SPI_ALT is

	signal RX_32BIT_SREG, N_RX_32BIT_SREG 			: STD_LOGIC_VECTOR(31 DOWNTO 0);		-- 32 BIT SHIFT REGISTER DEDICATED FOR ACTIVE SPI RECEIVE
	
	attribute syn_preserve : boolean;
	attribute syn_preserve of RX_32BIT_SREG : signal is true;
	attribute syn_preserve of N_RX_32BIT_SREG : signal is true;

	signal TX_32BIT_SREG, N_TX_32BIT_SREG 			: STD_LOGIC_VECTOR(31 DOWNTO 0);		-- 32 BIT SHIFT REGISTER DEDICATED FOR ACTIVE SPI TRANSMIT
	
	SIGNAL TX_32BIT_REG, N_TX_32BIT_REG				: STD_LOGIC_VECTOR(31 DOWNTO 0);		-- 32 BIT FIXED REGISTER DEDICATED FOR ACTIVE SPI TRANSMIT
	
	SIGNAL CLK_FCNT, N_CLK_FCNT						: INTEGER RANGE 0 TO 32;				-- SPI FRAME COUNTER
	SIGNAL CLK_FCNT_1C, CLK_FCNT_2C					: INTEGER RANGE 0 TO 32;				-- USED FOR CLOCK BOUNDARY CROSSING
	
	SIGNAL I_SCA_DAT_IN, N_I_SCA_DAT_IN				: STD_LOGIC;							-- INTERNAL SIGNAL FOR SCA TX SERIAL DATA LINE
	
	SIGNAL SPI_CLR, N_SPI_CLR						: STD_LOGIC;							-- SIGNAL USED TO CLEAR SPI REGSITERS
	SIGNAL CLK_FCNT_EN, N_CLK_FCNT_EN				: STD_LOGIC;							-- ENABLE FOR THE FRAME COUNTER
	SIGNAL I_SPI_RX_STRB, N_I_SPI_RX_STRB 			: STD_LOGIC;							-- SINGLE CLOCK PULSE STROBE INDICATES NEW SPI WORD RECEIVED
	SIGNAL I_SPI_RX_WORD, N_I_SPI_RX_WORD 			: STD_LOGIC_VECTOR(31 DOWNTO 0);		-- INTERNAL 32 BIT SHIFT REGISTER DEDICATED FOR ACTIVE SPI RECEIVE
	
	-- DEFINE THE STATES FOR THE MACHINE STATE MANAGING THE SPI PORT
	TYPE SPI_SM_STATES IS (INIT, DET_NULLCLK, EN_DET_FRAME1CNT, PIPELINE_DELAY, DET_FRAME_DONE, PROCESS_FRAME);	
	SIGNAL SPI_SM, N_SPI_SM							: SPI_SM_STATES;
	
	SIGNAL SCA_CLK_OUT_1C, SCA_CLK_OUT_2C			: STD_LOGIC;							-- USED FOR CLOCK BOUNDARY CROSSING
	
	SIGNAL NULLCLK_CNT, N_NULLCLK_CNT 				: INTEGER RANGE 0 TO 31;				-- COUNT OF THE NUMBER OF CLK-NULL SAMPLES

-- FOR DEBUG	
	SIGNAL STATE_ID 								: STD_LOGIC_VECTOR(3 DOWNTO 0);
begin

-- architecture body

--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE THE SPI INPUT AND OUTPUT DATA SHIFT REGISTERS WHICH OPERATES DIRECTLY FROM THE SPI CLOCK
-- DEFINE THE FRAME COUNT WHICH COUNTS CLOCK CYCLES DURING THE ACTIVE CLOCK CYCLES OF A 32-CYCLE DATA FRAME
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE THE D FF'S
SREG_DFF:PROCESS(SCA_CLK_OUT, SPI_CLR)
	BEGIN
		IF SPI_CLR = '1' THEN																-- AN EXTERNAL STATE MACHINE FORCES SYNCHRONIZATION OF THE SPI 
			RX_32BIT_SREG							<=	(OTHERS => '0');
			TX_32BIT_SREG							<=	(OTHERS => '0');
			CLK_FCNT								<=	 0;									-- FIRST TRANSITION GOES TO 1
			
			I_SCA_DAT_IN							<=	'0';
			
		ELSIF RISING_EDGE(SCA_CLK_OUT) THEN
			RX_32BIT_SREG							<=	N_RX_32BIT_SREG;
			TX_32BIT_SREG							<=	N_TX_32BIT_SREG;
			CLK_FCNT								<=	N_CLK_FCNT;
			
			I_SCA_DAT_IN							<=	N_I_SCA_DAT_IN;
			
		END IF;
	
	END PROCESS;

-- DEFINE D FF INPUTS THAT OPERATE DIRECTLY OFF THE SPI CLOCK HERE
SREG_DFFI:PROCESS(RX_32BIT_SREG, SCA_DAT_OUT, CLK_FCNT, CLK_FCNT_EN, TX_32BIT_REG, TX_32BIT_SREG)
	BEGIN	
		-- THIS IS THE RX PATH
		N_RX_32BIT_SREG(31 DOWNTO 0)				<=	RX_32BIT_SREG(30 DOWNTO 0) & SCA_DAT_OUT;		-- THESE ARE THE D FF INPUTS FOR THE SHIFT REGISTER 
																										-- SCA SPI SENDS MSb FIRST TO THE FPGA

		-- THIS COUNTS THE FRAME BITS
		IF CLK_FCNT = 32 THEN
			N_CLK_FCNT		<=	0;															-- NORMAL COUNT OP IS 1 THRU 32,WHERE 0 IS A HOLD / INIT VAL
		ELSIF CLK_FCNT_EN = '1'		THEN													-- THIS COUNTS THE SERIAL FRAME CLOCK CYCLES WHEN ENABLED
			N_CLK_FCNT								<=	CLK_FCNT + 1;			
		ELSE
			N_CLK_FCNT								<=	CLK_FCNT;
		END IF;

		N_I_SCA_DAT_IN							<=	TX_32BIT_SREG(31);						-- FPGA SPI SENDS MSb OUT FIRST TO SCA
		
		N_TX_32BIT_SREG							<=	TX_32BIT_SREG;						-- DEFAULT ASSIGNMENT
		
		CASE CLK_FCNT IS
			WHEN 0 =>	
				N_TX_32BIT_SREG					<=	TX_32BIT_REG;						-- *** SAMPLE EXTERAL DATA TO BE TRANSMITTED HERE ***
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(31);					-- FPGA SPI SENDS MSb OUT FIRST TO SCA
			WHEN 1 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(30);
			WHEN 2 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(29);
			WHEN 3 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(28);
			WHEN 4 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(27);
			WHEN 5 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(26);
			WHEN 6 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(25);
			WHEN 7 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(24);
			WHEN 8 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(23);
			WHEN 9 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(22);
			WHEN 10 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(21);
			WHEN 11 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(20);
			WHEN 12 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(19);
			WHEN 13 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(18);
			WHEN 14 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(17);
			WHEN 15 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(16);
			WHEN 16 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(15);
			WHEN 17 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(14);
			WHEN 18 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(13);
			WHEN 19 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(12);
			WHEN 20 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(11);
			WHEN 21 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(10);
			WHEN 22 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(9);
			WHEN 23 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(8);
			WHEN 24 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(7);
			WHEN 25 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(6);
			WHEN 26 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(5);
			WHEN 27 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(4);
			WHEN 28 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(3);
			WHEN 29 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(2);
			WHEN 30 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(1);
			WHEN 31 =>	
				N_I_SCA_DAT_IN					<=	TX_32BIT_SREG(0);
				
		END CASE;

		

	END PROCESS;


--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE THE REGISTERS THAT OPERATE FROM THE 5 MHZ CLOCK

REG_5M:PROCESS(CLK5M_OSC, MASTER_RST_B)
		BEGIN
			
			IF MASTER_RST_B = '0'  THEN
				SPI_SM				<=	INIT;
				CLK_FCNT_EN			<=	'0';
				SPI_CLR				<=	'0';
				I_SPI_RX_STRB		<=	'0';
				I_SPI_RX_WORD		<=	(OTHERS => '0');

				CLK_FCNT_1C			<=	 0;
				CLK_FCNT_2C			<=   0;
				
				SCA_CLK_OUT_1C		<=	'0';
				SCA_CLK_OUT_2C		<=	'0';
				
				NULLCLK_CNT			<=	 0;
				
				TX_32BIT_REG		<=	(OTHERS => '0');

			ELSIF RISING_EDGE(CLK5M_OSC)	THEN
				SPI_SM				<=	N_SPI_SM;
				CLK_FCNT_EN			<=	N_CLK_FCNT_EN;
				SPI_CLR				<=	N_SPI_CLR;
				I_SPI_RX_STRB		<=	N_I_SPI_RX_STRB;
				I_SPI_RX_WORD		<=	N_I_SPI_RX_WORD;

				CLK_FCNT_1C			<=	CLK_FCNT;						-- CLOCK BOUNDARY CROSSING
				CLK_FCNT_2C			<=	CLK_FCNT_1C;					-- CLOCK BOUNDARY CROSSING
				
				SCA_CLK_OUT_1C		<=	SCA_CLK_OUT;					-- CLOCK BOUNDARY CROSSING
				SCA_CLK_OUT_2C		<=	SCA_CLK_OUT_1C;					-- CLOCK BOUNDARY CROSSING
				
				NULLCLK_CNT			<=	N_NULLCLK_CNT;
				
				TX_32BIT_REG		<=	N_TX_32BIT_REG;
			
			END IF;
END PROCESS;


--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--  THIS PROCESS CONTROLS THE SPI INPUT AND OUTPUT SHIFT REGISTERS AS WELL AS THE SPI CLOCK COUNT FOR THE FRAME
--  CLOCK BOUNDARY CROSSING IS INHERENTLY SYNCHRONOUS FOR THE CONTROL SIGNALS ONCE THE STATE MACHINE IS SYNCHRONIZED TO THE SPI FRAME
--  HOWEVER, DOUBLE REGISTERS ARE USED TO SAMPLE THE CLK_FCNT AS WELL AS THE SPI CLOCK

SPI:PROCESS(SPI_SM, CLK_FCNT_2C, SCA_CLK_OUT_2C, RX_32BIT_SREG, NULLCLK_CNT, I_SPI_RX_WORD, CLK_FCNT_EN, SPI_CLR, SPI_TX_WORD, TX_32BIT_REG,
			STATE_ID)
	BEGIN
	
		-- DEFAULT ASSIGNMENTS THAT GET OVER-WRITTEN BELOW AS NEEDED:
		N_NULLCLK_CNT		<=	NULLCLK_CNT;
		N_I_SPI_RX_STRB		<=	'0';
		N_SPI_CLR			<=	SPI_CLR;
		N_CLK_FCNT_EN		<=	CLK_FCNT_EN;
		N_I_SPI_RX_WORD		<=  I_SPI_RX_WORD;
		N_TX_32BIT_REG		<=	TX_32BIT_REG;

		CASE SPI_SM IS
	
			WHEN INIT	=>

				N_CLK_FCNT_EN		<=	'0';						-- DISABLE TO THE FRAME COUNTER
				N_SPI_CLR			<=	'1';						-- SEND OUT A CLEAR TO INITIALIZE THE FRAME COUNTER AND SPI INPUT DATA REGISTER

				N_SPI_SM			<=	DET_NULLCLK; 				-- GO WAIT FOR DETECTION OF A NULL CLOCK CONDITION TO SYNCH THE SPI FRAME

				N_NULLCLK_CNT		<=	0;							-- INITIALIZE THE NULL CLOCK COUNTER
				
				STATE_ID	<=	"0000";
		
			WHEN DET_NULLCLK	=>									-- WAIT HERE UNTIL THE SPI CLOCK IS NULL FOR AT LEASTY 3/4 SPI CLOCK PERIOD
				N_CLK_FCNT_EN		<=	'0';						-- DISABLE TO THE FRAME COUNTER
				N_SPI_CLR			<=	'1';						-- SEND OUT A CLEAR TO INITIALIZE THE FRAME COUNTER AND SPI INPUT DATA REGISTER
				
				IF NULLCLK_CNT > 17	THEN							-- ONE SPI CLOCK PERIOD COUNT WHILE HIGH IS 5MHZ/312KHZ/2 = ~ 8 COUNTS
					N_NULLCLK_CNT		<=	0;						-- IF NULL CLOCK, THEN CLEAR THE CNT
					N_SPI_SM			<=	EN_DET_FRAME1CNT;		-- AND GO WAIT FOR THE NEXT FRAME TO BE COMPLETED

				ELSIF	SCA_CLK_OUT_2C = '0'	THEN				-- ONLY COUNT DURING THE LOGIC LOW PORTION OF THE SPI CLOCK SIGNAL
					N_NULLCLK_CNT		<=  NULLCLK_CNT + 1;
					N_SPI_SM			<=	DET_NULLCLK;			-- STAY HERE UNTIL NULL DETECTED
					
				ELSE
					N_NULLCLK_CNT		<=	0;						-- ONLY GET HERE IF THE SPI CLOCK IS ACTIVE
					N_SPI_SM			<=	DET_NULLCLK;			-- STAY HERE UNTIL NULL DETECTED
					
				END IF;
				
				STATE_ID	<=	"0001";

		 
			WHEN EN_DET_FRAME1CNT	=>								-- ENABLE THE DET FRAME CNT AND ALSO RELEASE THE CLEAR
				N_CLK_FCNT_EN		<=	'1';						-- ENABLE THE FRAME COUNTER
				N_SPI_CLR			<=	'0';						-- DISABLE THE SPI_CLR
				N_SPI_SM			<=	PIPELINE_DELAY;				-- GO WAIT ONE MORE CLOCK CYCLE TO ALLOW FOR THE CLOCK BOUNDARY CROSSING
			
				STATE_ID	<=	"0010";

			
			WHEN PIPELINE_DELAY	=>									-- NEED A PIPELINE DELAY TO ACCOUNT FOR THE CLOCK BOUNDARY CROSSING REGISTERS
				N_SPI_SM			<=	DET_FRAME_DONE;
				
				STATE_ID	<=	"0011";
			
			WHEN DET_FRAME_DONE =>									-- WAIT HERE UNTIL 32 SPI CLOCK PERIODS HAVE BEEN DETECTED.
		 
	
				IF CLK_FCNT_2C	=  32	THEN
					N_SPI_SM			<=	PROCESS_FRAME;
				ELSE
					N_SPI_SM			<=	DET_FRAME_DONE;
				END IF;
				
				N_TX_32BIT_REG		<=	SPI_TX_WORD;				-- COPY THE DATA WORD TO BE TRANSMITTED DURING NEXT FRAME INTO A REGISTER
				
				STATE_ID	<=	"0100";
				
			WHEN PROCESS_FRAME	=>	
				N_I_SPI_RX_WORD		<= RX_32BIT_SREG;				-- SEND OUT A COPY THE RECEIVED SERIAL 32 BIT WORD
				N_I_SPI_RX_STRB		<=	'1';						-- SINGLE CLOCK PULSE STROBE INDICATES NEW FRAME READY
				N_SPI_SM			<=	INIT;
			
				STATE_ID	<=	"0101";
				
			
			WHEN OTHERS			=>
				N_SPI_SM			<=	INIT;
			
				STATE_ID	<=	"0110";
				
		END CASE;

	END PROCESS;
	
-- ASSIGN INTERNAL SIGNALS TO EXTERNAL PORTS
SPI_RX_STRB		<=	I_SPI_RX_STRB;
SPI_RX_WORD		<=	I_SPI_RX_WORD;

SCA_DAT_IN		<=	I_SCA_DAT_IN;
P_STATE_ID		<=	STATE_ID;

P_TX_32BIT_REG	<=	TX_32BIT_REG;

end RTL;
