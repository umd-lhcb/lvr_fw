--------------------------------------------------------------------------------
-- Company: UNIVERSITY OF MARYLAND
--
-- File: SERIAL_RX.vhd
-- File history:
--      <Rev - // Mar 28, 2017  INITIAL
--
-- Description: THIS MODULE RECEIVES THE SERIAL WORD.
--					FRAME PACKET CONSISTS OF 16 BITS + 2 START AND 2 STOP BITS.
--					LSB ASSUMED FIRST
--					THE START AND STOP BITS ARE ALL LOGIC '1'
--					15		ODD PARITY (APPLIES TO DATA BITS ONLY)
--					14		UVL STATUS
--					13..12	MODE 
--					11..8	MODULE ADDRESS
--					7..0	CHANNEL ENABLES
--					
--					
--					BIT IS DERIVED FROM 5 MHZ CLOCK DIVIDED BY 64 = 12.8 USEC (78.125 KBPS)
--					12.8 USEC / 200NS = 64 COUNTS
--
--					THE RX_INPUT IS ASSUMED TO BE DIGITALLY FILTERED TO ELIMINATE ANY SPIKES/GLITCHES/ETC.....
--
-- Targeted device: <Family::ProASIC3> <Die::A3PN125> <Package::100 VQFP>
-- Author: TOM O'BANNON
--
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_MISC.ALL;
USE IEEE.NUMERIC_STD.ALL;

library proasic3;
use proasic3.all;

-- NOTE:  THE SYNPLIFY LIBRARY NEEDS TO BE COMMENTED OUT FOR MODELSIM PRESYNTH SIMS SINCE MODELSIM DOES NOT RECOGNIZE IT
library synplify;
use synplify.attributes.all;

entity SERIAL_RX is
port (
		MASTER_RST_B		:	IN	STD_LOGIC;							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
		CLK_5M_GL			:	IN	STD_LOGIC;
		RX_INPUT			:	IN	STD_LOGIC;							-- FINAL RX SIGNAL BIT STREAM AFTER THE FILTER FUNCTION AND HYSTERISIS HAVE BEEN APPLIED
		MODULE_ADDR			:	IN	STD_LOGIC_VECTOR(4 DOWNTO 0);		-- HARDWIRED ADDRESS OF THIS MODULE
		
		RX_WORD				:	OUT	STD_LOGIC_VECTOR(14 DOWNTO 0);		-- FINAL RECEIVED RX WORD (BIT 15 IN RX BIT STREAM IS PARITY PLACEHOLDER)
		RX_ODD_PARITY		:	OUT	STD_LOGIC;							-- ODD PARITY FOR THE RX_WORD (FOR SIM DEBUG)
		RX_PARITY_ERR		:	OUT	STD_LOGIC;							-- LATCHED VESRION OF THE LAST RX PARITY ERROR
		RX_STRB				:	OUT	STD_LOGIC							-- SINGLE CLOCK PULSE STRB INDICATES THE RX_WORD WAS UPDATED AND HAS NO PARITY ERROR
	);
end SERIAL_RX;

architecture RTL of SERIAL_RX is
ATTRIBUTE SYN_RADHARDLEVEL OF RTL : ARCHITECTURE IS "TMR";

-- !!!!!  NOTE   !!!! THE STATE MACHINES NEED TO HAVE THE "SAFE ATTRIBUTE" APPLIED IN SYNTHESIS

-- DEFINE THE STATES FOR SERIAL RECEIVE STATE MACHINE-----!!!!! ADD PLACEHOLDERS TO CREATE 2^^N STATES !!!!!!
TYPE RECEIVE_STATES IS (	INIT, BIT_DEL_WAIT, DET_1ST_START_BIT, DET_2ND_START_BIT, 
					RX_0LS_BIT, RX_1_BIT, RX_2_BIT, RX_3_BIT, RX_4_BIT, RX_5_BIT, RX_6_BIT, RX_7_BIT, 
					RX_8_BIT, RX_9_BIT, RX_10_BIT, RX_11_BIT, RX_12_BIT, RX_13_BIT, RX_14_BIT, RX_15_BIT, 
					DET_1ST_STOP_BIT, DET_2ND_STOP_BIT, CHECK_PARITY, CHECK_M_ADDR, FINISH_STROBE
					);

SIGNAL 	N_RX_STATE, RX_STATE 				: 	RECEIVE_STATES;								-- STATE MACHINE COUNTER FOR THE RX STATE MACHINE
SIGNAL	N_RET_STATE, RET_STATE				:	RECEIVE_STATES;								-- POINTER FOR A RETURN LOCATION ON THE RX STATE MACHINE

SIGNAL	N_BIT_POSN_CNT, BIT_POSN_CNT		:	INTEGER RANGE 0 TO 127;						-- COUNTER USED TO MEASURE BIT POSITION EVENTS
SIGNAL	N_SER_WORD, SER_WORD				:	STD_LOGIC_VECTOR(15 DOWNTO 0);				-- RECEIVED SERIAL WORD BUFFER
SIGNAL	N_WORD_STRB, WORD_STRB				:	STD_LOGIC;									-- STROBE PULSE, 1 CLOCK WIDE, INDICATES NEW RX WORD READY
SIGNAL	N_ODD_PARITY, ODD_PARITY			:	STD_LOGIC;									-- ODD PARITY BIT FOR RX WORD

SIGNAL 	N_PARITY_ERR, PARITY_ERR			:	STD_LOGIC;									-- LATCHED VERSION OF LAST RX PARITY ERROR CONDITION

CONSTANT	HALF_BIT_CNT					:	INTEGER RANGE 0 TO 127 := 29;				-- 32 COUNTS OF 5 MHZ CLOCK = 1/2 SERIAL BIT POSITION
CONSTANT 	FULL_BIT_CNT					:	INTEGER RANGE 0 TO 127 := 61;				-- 64 COUNTS OF 5 MHZ CLOCK = FULL SERIAL BIT POSITION

begin

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE ALL REGISTERS USED WITH THE 5 MHZ CLOCK
REG5M:PROCESS(CLK_5M_GL, MASTER_RST_B)	
	BEGIN
		IF MASTER_RST_B = '0' THEN
			RX_STATE		<=	INIT;
			BIT_POSN_CNT	<=	 0;
			SER_WORD		<=	(OTHERS => '0');
			WORD_STRB		<=	'0';
			ODD_PARITY		<=	'0';
			PARITY_ERR		<=	'0';
			RET_STATE		<=	INIT;
			
		ELSIF (CLK_5M_GL'EVENT AND CLK_5M_GL='1') THEN
			RX_STATE		<=	N_RX_STATE;
			BIT_POSN_CNT	<=	N_BIT_POSN_CNT;
			SER_WORD		<=	N_SER_WORD;
			WORD_STRB		<=	N_WORD_STRB;
			ODD_PARITY		<=	N_ODD_PARITY;
			PARITY_ERR		<=	N_PARITY_ERR;
			RET_STATE		<=	N_RET_STATE;
			
		END IF;
		
	END PROCESS;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE THE SERIAL RX PROCESS
SER_RX:PROCESS(RX_STATE, RET_STATE, BIT_POSN_CNT, RX_INPUT, SER_WORD, ODD_PARITY, WORD_STRB, MODULE_ADDR, PARITY_ERR)
	BEGIN
	
	-- DEFAULT ASSIGNMENTS (GET OVER-WRITTEN BELOW AS NEEDED)
	N_RET_STATE			<=	RET_STATE;
	N_BIT_POSN_CNT		<=	BIT_POSN_CNT;
	N_ODD_PARITY		<=	ODD_PARITY;
	N_SER_WORD			<=	SER_WORD;
	N_WORD_STRB			<=	WORD_STRB;
	N_PARITY_ERR		<=	PARITY_ERR;
	
		CASE RX_STATE IS

			WHEN INIT			=>								-- WAIT HERE FOR A LOGIC 1 DETECTION ON THE RX_INPUT
				IF RX_INPUT = '1'	THEN
					N_RX_STATE		<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
					N_RET_STATE		<=	DET_1ST_START_BIT;		-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
					N_BIT_POSN_CNT	<=	HALF_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE HALF BIT COUNT VALUE
				ELSE
					N_RX_STATE		<=	INIT;					-- STAY HERE UNLESS '1' DETECTED ON RX_INPUT
					N_RET_STATE		<=	INIT;					-- INITIALIZE THE POINTER TO THE RETURN STATE WHEN COUNTING BIT DELAYS
					N_BIT_POSN_CNT	<=	BIT_POSN_CNT;
				END IF;

				N_ODD_PARITY	<=	 '0';						-- INITIALIZE THE RX ODD PARITY BIT

			WHEN BIT_DEL_WAIT	=>								-- WAIT HERE FOR THE SPECIFIED BIT TIME DELAY--THIS STATE STEP IS REUSED TO MEASURE EACH 1 OR 1/2 BIT DURATION
				IF  BIT_POSN_CNT = 0	THEN
					N_RX_STATE		<=	RET_STATE;				-- BRANCH TO THE NEXT STATE
					N_RET_STATE		<=	RET_STATE;				-- JUST STORE CURRENT VALUE
					N_BIT_POSN_CNT	<=	BIT_POSN_CNT;			-- JUST STORE CURRENT VALUE
				ELSE
					N_RX_STATE		<=	BIT_DEL_WAIT;			-- STAY HERE UNTIL DONE
					N_RET_STATE		<=	RET_STATE;				-- JUST STORE CURRENT VALUE
					N_BIT_POSN_CNT	<=	BIT_POSN_CNT - 1;		-- DECREMENT THE COUNTER
				END IF;
				
			WHEN DET_1ST_START_BIT	=>							-- TEST FOR THE FIRST START BIT
				IF RX_INPUT = '1'	THEN
					N_RX_STATE		<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
					N_RET_STATE		<=	DET_2ND_START_BIT;		-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
					N_BIT_POSN_CNT	<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				ELSE
					N_RX_STATE		<=	INIT;					-- GO BACK TO INIT IF A '1' IS NOT DETECTED ON THE RX_INPUT
					N_RET_STATE		<=	INIT;					-- INITIALIZE THE POINTER TO THE RETURN STATE WHEN COUNTING BIT DELAYS
					N_BIT_POSN_CNT	<=	BIT_POSN_CNT;			-- JUST STORE CURRENT VALUE
				END IF;
				
			WHEN DET_2ND_START_BIT	=>							-- TEST FOR THE SECOND START BIT
				IF RX_INPUT = '1'	THEN						-- IF THERE, THEN STORE THE NEXT 16 DATA BITS
					N_RX_STATE		<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
					N_RET_STATE		<=	RX_0LS_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
					N_BIT_POSN_CNT	<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				ELSE
					N_RX_STATE		<=	INIT;					-- GO BACK TO INIT IF A '1' IS NOT DETECTED ON THE RX_INPUT
					N_RET_STATE		<=	INIT;					-- INITIALIZE THE POINTER TO THE RETURN STATE WHEN COUNTING BIT DELAYS
					N_BIT_POSN_CNT	<=	BIT_POSN_CNT;			-- JUST STORE CURRENT VALUE
				END IF;

			WHEN RX_0LS_BIT		=>								-- STORE THE LSB 0 BIT VALUE
				N_SER_WORD(0)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_1_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_1_BIT		=>								-- STORE THE LSB 1 BIT VALUE
				N_SER_WORD(1)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_2_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_2_BIT		=>								-- STORE THE LSB 2 BIT VALUE
				N_SER_WORD(2)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_3_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_3_BIT		=>								-- STORE THE LSB 3 BIT VALUE
				N_SER_WORD(3)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_4_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_4_BIT		=>								-- STORE THE LSB 4 BIT VALUE
				N_SER_WORD(4)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_5_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_5_BIT		=>								-- STORE THE LSB 5 BIT VALUE
				N_SER_WORD(5)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_6_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE

			WHEN RX_6_BIT		=>								-- STORE THE LSB 6 BIT VALUE
				N_SER_WORD(6)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_7_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_7_BIT		=>								-- STORE THE LSB 7 BIT VALUE
				N_SER_WORD(7)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_8_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_8_BIT		=>								-- STORE THE LSB 8 BIT VALUE
				N_SER_WORD(8)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_9_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_9_BIT		=>								-- STORE THE LSB 9 BIT VALUE
				N_SER_WORD(9)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_10_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_10_BIT		=>								-- STORE THE LSB 10 BIT VALUE
				N_SER_WORD(10)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_11_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_11_BIT		=>								-- STORE THE LSB 11 BIT VALUE
				N_SER_WORD(11)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_12_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_12_BIT		=>								-- STORE THE LSB 12 BIT VALUE
				N_SER_WORD(12)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_13_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_13_BIT		=>								-- STORE THE LSB 13 BIT VALUE
				N_SER_WORD(13)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_14_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_14_BIT		=>								-- STORE THE LSB 14 BIT VALUE
				N_SER_WORD(14)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	RX_15_BIT;				-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY XOR RX_INPUT;-- CALCULATE THE RUNNING PARITY

			WHEN RX_15_BIT		=>								-- STORE THE LSB 15 BIT VALUE---THIS IS THE PARITY BIT-- SO NO PARITY CALC NEEDED!!!!
				N_SER_WORD(15)		<=	RX_INPUT;
				N_RX_STATE			<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
				N_RET_STATE			<=	DET_1ST_STOP_BIT;		-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
				N_BIT_POSN_CNT		<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				N_ODD_PARITY		<=	ODD_PARITY ;			-- CALCULATE THE RUNNING PARITY
				

			WHEN DET_1ST_STOP_BIT	=>							-- TEST FOR THE FIRST STOP BIT
				IF RX_INPUT = '1'	THEN
					N_RX_STATE		<=	BIT_DEL_WAIT;			-- NEXT STATE IS TO COUNT THE SPECIFIED BIT POSITION TIME
					N_RET_STATE		<=	DET_2ND_STOP_BIT;		-- INITIALIZE THE POINTER TO THE NEXT RETURN STATE WHEN COUNTING BIT DELAYS
					N_BIT_POSN_CNT	<=	FULL_BIT_CNT;			-- INTIALIZE THE BIT SAMPLE POSITION COUNTER WITH THE FULL BIT COUNT VALUE
				ELSE
					N_RX_STATE		<=	INIT;					-- GO BACK TO INIT IF A '1' IS NOT DETECTED ON THE RX_INPUT
					N_RET_STATE		<=	INIT;					-- INITIALIZE THE POINTER TO THE RETURN STATE WHEN COUNTING BIT DELAYS
					N_BIT_POSN_CNT	<=	BIT_POSN_CNT;			-- JUST STORE CURRENT VALUE
				END IF;
				
			WHEN DET_2ND_STOP_BIT	=>							-- TEST FOR THE SECOND STOP BIT
				IF RX_INPUT = '1'	THEN						-- IF THERE, THEN GO CHECK THE PARITY
					N_RX_STATE		<=	CHECK_PARITY;			-- 
					N_RET_STATE		<=	RET_STATE;				-- JUST STORE CURRENT VALUE
					N_BIT_POSN_CNT	<=	BIT_POSN_CNT;			-- JUST STORE CURRENT VALUE
				ELSE
					N_RX_STATE		<=	INIT;					-- GO BACK TO INIT IF A '1' IS NOT DETECTED ON THE RX_INPUT
					N_RET_STATE		<=	INIT;					-- INITIALIZE THE POINTER TO THE RETURN STATE WHEN COUNTING BIT DELAYS
					N_BIT_POSN_CNT	<=	BIT_POSN_CNT;			-- JUST STORE CURRENT VALUE
				END IF;

			WHEN CHECK_PARITY		=>							-- LAST STEP IS TO CHECK THE PARITY BEFORE GENERATING A STROBE PULSE FOR THE NEW WORD
				IF ODD_PARITY	= SER_WORD(15)	THEN
					N_RX_STATE		<=	FINISH_STROBE;
					N_WORD_STRB		<=	'1';
					N_PARITY_ERR	<=	'0';
				ELSE
					N_RX_STATE		<=	INIT;					-- PARITY ERROR, THEREFORE IGNORE RX (FOR NOW)
					N_WORD_STRB		<=	'0';
					N_PARITY_ERR	<=	'1';
				END IF;
				
			WHEN CHECK_M_ADDR		=>							-- LAST STEP IS TO CHECK THE MODULE ADDRESS BEFORE GENERATING A STROBE PULSE FOR THE NEW WORD
				IF MODULE_ADDR	= SER_WORD(11 DOWNTO 8)	THEN
					N_RX_STATE		<=	FINISH_STROBE;
					N_WORD_STRB		<=	'1';
				ELSE
					N_RX_STATE		<=	INIT;					-- NOT THIS MODULE'S ADDR, THEREFORE IGNORE RX
					N_WORD_STRB		<=	'0';
				END IF;

			WHEN FINISH_STROBE		=>	
					N_RX_STATE		<=	INIT;					-- 
					N_WORD_STRB		<=	'0';
						
		END CASE;

	END PROCESS;
-- ASSIGN INTERNAL SIGNALS TO EXTERNAL PORTS 
RX_STRB			<=	WORD_STRB;
RX_WORD			<=	SER_WORD(14 DOWNTO 0);						-- BIT 15 IS PARITY
RX_ODD_PARITY	<=	ODD_PARITY;
RX_PARITY_ERR	<=	PARITY_ERR;
	
	
end RTL;
