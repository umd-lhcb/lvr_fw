--------------------------------------------------------------------------------
-- Company: UNIVERSITY OF MARYLAND
--
-- File: TOP_LV_REGUL_CNTL.vhd
-- File history:
--      REV - // JAN 7, 2019  INITIAL UPDATE
--
-- Description: LV REGULATOR SERIAL CONTROL INTERFACE
--      FUNCTIONS:
--          		1) UNDER-VOLTAGE LOCKOUT FAILSAFE--CHECK EACH OF 4 FUSES
--					2) BOARD OVER-TEMPERATURE FAILSAFE CHECK
--          		3) SERIAL COMM
--          		4) REGULATOR CHANNEL SEQUENCE CONTROLS

-- 		THERE ARE 2 SERIAL COMM OPTIONS:
--			(A) SINGLE GBT-SCA SPI SLAVE WHEN ADDR_SEL(4:0)= 1F HEX
--					NOTE THAT THIS SPI PORT OPERATES AS A SHIFT REGISTER DRIVEN BY THE GBT-SCA SPI CLOCK.  
--					A CLOCK BOUNDARY CROSSING IS INITIATED ONCE THE SPI CLOCK STOPS

--			(B) DAISY CHAINED RS-485 ASYNC SERIAL INTERFACE

--
-- Targeted device: <Family::ProASIC3N> <Die::A3PN250> <Package::100 VQFP>
-- Author: TOM O'BANNON
--
-- ////////////////////////////////////////////////////////////////////////////////////
-- ////////////////////////////////////////////////////////////////////////////////////
-- CAUTION:  SIM_MODE CONSTANT NEEDS TO BE MANUALLY UPDATED!!!!!
-- 				(A) SLOW_PULSE_EN_GEN HAS A SPECIAL SIM INPUT OPTION
--				(B) MAIN_SEQUENCER CONSTANT DEL_CNT_VAL CAN BE CHANGED TO SPPED SIM
-- ////////////////////////////////////////////////////////////////////////////////////
-- ////////////////////////////////////////////////////////////////////////////////////
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_MISC.ALL;
--USE IEEE.NUMERIC_STD.ALL;

library proasic3;
use proasic3.all;

-- NOTE:  THE SYNPLIFY LIBRARY NEEDS TO BE COMMENTED OUT FOR MODELSIM PRESYNTH SIMS SINCE MODELSIM DOES NOT RECOGNIZE IT
library synplify;
use synplify.attributes.all;

entity TOP_LV_REGUL_CNTL is
port (
        CLK40M_OSC          	:   IN  STD_LOGIC;                      	-- pin 57, EXTERNAL 3.3V 40 MHZ CLOCK 
        POR_FPGA            	:   IN  STD_LOGIC;                         	-- pin 93, ACTIVE LOW RESET --DEDICATED RC TIME CONSTANT---NEEDS SCHMITT-TRIGGER!

-- UNDER-VOLTAGE LOCKOUT AND FUSE STATUS DETECTION	
		FPGA_FUSE_1_2_OK		:	IN	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- pin 42, UNDER-VOLTAGE LOCKOUT FAILSAFE INPUT ('1'= INPUT FUSED RAIL FOR CH1&2 ABOVE THRESHOLD)
		FPGA_FUSE_3_4_OK		:	IN	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- pin 41, UNDER-VOLTAGE LOCKOUT FAILSAFE INPUT ('1'= INPUT FUSED RAIL FOR CH3&4 ABOVE THRESHOLD)
		FPGA_FUSE_5_6_OK		:	IN	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- pin 40, UNDER-VOLTAGE LOCKOUT FAILSAFE INPUT ('1'= INPUT FUSED RAIL FOR CH5&6 ABOVE THRESHOLD)
		FPGA_FUSE_7_8_OK		:	IN	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- pin 36, UNDER-VOLTAGE LOCKOUT FAILSAFE INPUT ('1'= INPUT FUSED RAIL FOR CH7&8 ABOVE THRESHOLD)

-- OVER-TEMPERATURE FAILSAFE
		TEMP_OK_B				:	IN	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- pin 43, BOARD TEMPERATURE FAILSAFE OK ('0'= ABOVE THE OVER-TEMP THRESHOLD)

-- DIP SWITCH INPUTS
	
	-- OPERATION AND FAILSAFE MODES: DIP SW SETTINGS
		MODE_2					:	IN	STD_LOGIC;							-- pin 31, OP MODE			'1' = SPECIAL TEST LOW DUTY CYCLE MODE
																			--   						'0' = NORMAL OP WITH STAGGERED ENABLE SEQUENCES (19.6608 MS PER CHANNEL)
		MODE_1					:	IN	STD_LOGIC;							-- pin 30, WDT_EN			'1' = WATCH DOG TIMER ENABLED
																			--	 						'0' = WATCH DOG TIMER DISABLED
		MODE_0					:	IN	STD_LOGIC;							-- pin 29, DIAGNOSTIC MODE	'1' = DISABLE FRAME ERROR CHECKING
																			--							'0' = NORMAL OPERATION FRAME ERROR CHECK ENABLED
	-- MASTER-SLAVE CHANNEL GROUP ENABLES: DIP SW SETTINGS
	-- '0' = DISABLED STATE WHERE SPECIFIED CHANNELS TREATED INDEPENDENTLY	
	-- '1' = ENABLED STATE WHERE SPECIFIED CHANNELS ARE TREATED AS A MASTER-SLAVE PAIR	
		CH1_2_MS_CFG_EN			:	IN	STD_LOGIC;							-- pin 21, BIT 0:	CH1_2_MS_CFG_EN = CHANNELS 1 & 2
		CH3_4_MS_CFG_EN			:	IN	STD_LOGIC;							-- pin 20, BIT 1:	CH3_4_MS_CFG_EN = CHANNELS 3 & 4
		CH5_6_MS_CFG_EN			:	IN	STD_LOGIC;							-- pin 19, BIT 2:	CH5_6_MS_CFG_EN = CHANNELS 5 & 6
		CH7_8_MS_CFG_EN			:	IN	STD_LOGIC;							-- pin 16, BIT 3:	CH7_8_MS_CFG_EN = CHANNELS 7 & 8

	-- MANUAL CHANNEL GROUP ENABLES FOR STAND-ALONE TESTS:  DIP SW SETTINGS
		MAN_EN_CH_4TO1			:	IN	STD_LOGIC;							-- pin 15, (Schema was CH5_6_W_STDBY_E) NCHANNELS 5 & 6 TREATED AS REDUNDANT PAIR WHNE ='1'
		MAN_EN_CH_8TO5			:	IN	STD_LOGIC;							-- pin 13, (Schema was CH7_8_W_STDBY_EN) CHANNELS 7 & 8 TREATED AS REDUNDANT PAIR WHNE ='1'

		TEMP_FAILSAFE_EN		:	IN	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- pin 11, '1' = TEMPERATURE FAILSAFE IS ENABLED
		STDBY_OP_B				:	IN	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- PIN 10, '0'=NORMAL OP, '1'= FORCED V_OS OUT (was UVL_FAILSAFE_EN) '1' = UNDER-VOLTAGE LOCKOUTS ARE ENABLED (SPECIFIES THE MIN VOLTAGE REQUIRED TO OPERATE CHANNELS
	
-- RS-485		
		RX_FPGA					:	IN	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- pin 97, RS_485 SERIAL RX STREAM
		TX_FPGA					:	OUT	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- pin 98, RS_485 SERIAL TX STREAM
		
		PRI_RX_EN_BAR			:	OUT	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- pin 96, ENABLE FOR THE RX OUTPUT--SHOULD BE STUCK AT '0'
		PRI_TX_EN				:	OUT	STD_LOGIC;							-- pin 94, ENABLE FOR THE TX OUTPUT--
		
		ADDR_SEL			    :	IN	STD_LOGIC_VECTOR(4 DOWNTO 0);		-- pins {28, 27, 26, 23, 22} DIP SW FOR MODULE ADDRESS--THIS IS ONLY NEEDED FOR THE DAISY-CHAINED RS-485 INTERFACE

-- GBT-SCA SPI
		SCA_CLK_OUT				:	IN	STD_LOGIC;							-- pin 35, SPI CLOCK FROM THE SPI MASTER
		SCA_RESET_OUT			:	IN	STD_LOGIC;							-- pin 34, OPTIONAL RESET FROM THE SPI MASTER
		SCA_DAT_IN				:	OUT	STD_LOGIC;							-- pin 3, SERIAL DATA FROM FPGA TO THE SPI MASTER
		SCA_DAT_OUT				:	IN	STD_LOGIC;							-- pin 2, SERIAL DATA TO THE FPGA FROM THE SPI MASTER
		POR_OUT_TO_SCA			:	OUT	STD_LOGIC;							-- pin 6, RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE

		
-- CHANNEL ENABLES
		P_CH_MREG_EN			:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);		-- pins {62, 65, 71, 76, 80, 83, 92, 86} CHANNEL ENABLE SIGNAL: MAIN REGULATOR IC, ACTIVE HIGH
		P_CH_IAUX_EN			:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);		-- pins {61, 64, 70, 73, 79, 82, 85, 90} CHANNEL ENABLE SIGNAL: IAUX REGULATOR IC, ACTIVE HIGH
		P_CH_VOSG_EN			:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);		-- pins {60, 63, 69, 72, 78, 81, 84, 91} CHANNEL ENABLE SIGNAL: VOS_GEN REGULATOR IC, ACTIVE HIGH

-- MONITOR AND STATUS SIGNALS
		PWR_OK_LED				:	OUT	STD_LOGIC;							-- pin 95, 	STATUS YELLOW LED INDICATING AT LEAST ONE CHANNEL IS ACTIVE
																			-- 			SINGLE BLINK - CHANNEL ENABLE / DISABLE EVENT
		STATUS_LED				:	OUT	STD_LOGIC;							-- pin 77, 	STEADY=UVL'S OK, SINGLE BLINK=SEU AND/OR WDT

-- DIAGNOSTIC & TEST I/O
		BUF5M_J11_15_TCONN		:	OUT	STD_LOGIC;							-- PIN 35, (SCHEMA ALIAS= CS2_SEL_EN) 5 MHZ CLOCK BUFFER
		
-- UNUSED FPGA I/O BEING TIED TO SPECIFIED SAFE STATE
		UNUSED_1				:	IN	STD_LOGIC;							-- PIN 59, 3V3 BANK, NOT ROUTED FOR USE, BUT HAS 3V3 PULLUP PRESENT
		UNUSED_2				:	IN	STD_LOGIC;							-- PIN 58, 3V3 BANK, NOT ROUTED FOR USE, BUT HAS GND PULLDN PRESENT
		J11_25_TCONN			:	IN	STD_LOGIC;							-- pin 45, (SCHEMA ALIAS= SCLK_BUS)
		J11_27_TCONN			:	IN	STD_LOGIC;							-- pin 44, (SCHEMA ALIAS= SDAT_BUS)
		J11_17_TCONN			:	OUT	STD_LOGIC;							-- PIN 32, (SCHEMA ALIAS= CS3_SEL_EN) UNUSED I/O PIN
		J11_19_TCONN			:	OUT	STD_LOGIC;							-- PIN 8,  (SCHEMA ALIAS= CS4_SEL_EN) UNUSED I/O PIN
		J11_21_TCONN			:	OUT	STD_LOGIC;							-- PIN 7,  (SCHEMA ALIAS= CS5_SEL_EN) UNUSED I/O PIN
		J11_23_TCONN			:	OUT	STD_LOGIC							-- PIN 5,  (SCHEMA ALIAS= CS6_SEL_EN) UNUSED I/O PIN
        );

end TOP_LV_REGUL_CNTL;

architecture RTL of TOP_LV_REGUL_CNTL is


--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

-- ATTRIBUTE SYN_RADHARDLEVEL OF RTL : ARCHITECTURE IS "TMR";

--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++



--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- NOTES:  !!!!!	SPECIFIC I/O FEATURES (EG HYSTERISIS ) NEED TO BE ASSIGNED IN THE CONSTRAINTS FILE  !!!!
--		   !!!!!	THE SYN_ENCODING FOR EACH OF THE STATE MACHINES NEEDS TO HAVE A "SAFE, ORIGINAL" fsm ENCODING SEPECIFIED IN THE SYNTH CONSTRAINT FILE     !!!!!!!
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++


--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE COMPONENTS
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

-- IIR FILTER WITH SEVERAL USES:
-- 		(1) THE RS-485 SERIAL RECEIVE SIGNAL (ONLY--NOT USED FOR THE GBT-SCA SPI SLAVE PORT)		FILTERED RESULT:  FILTD_RS485RX
--		(2) TEMP_OK_B																				FILTERED RESULT:  FILTD_TEMP_OK_B
--		(3) FPGA_FUSE_X_Y_OK (4 FILTERS FOR 4 SIGNALS)												FILTERED RESULTS: FILTD_FUSE_X_Y_OK
COMPONENT IIR_FILT IS
port (
		MASTER_RST_B		:	IN	STD_LOGIC;							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
		CLK_5M_GL			:	IN	STD_LOGIC;
		
		SIG_IN				:	IN	STD_LOGIC_VECTOR(0 DOWNTO 0);		-- INPUT SIGNAL TO BE FILTERED
		THRESH_UPPER		:	IN	STD_LOGIC_VECTOR(7 DOWNTO 0);		-- UPPER HYSTERISIS THRESHOLD (IE RISING SIGNAL THRESHOLD)
		THRESH_LOWER		:	IN	STD_LOGIC_VECTOR(7 DOWNTO 0);		-- LOWER HYSTERISIS THRESHOLD (IE FALLING SIGNAL THRESHOLD)
		FILT_SIGOUT			:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);		-- RESULTING SIGNAL FILTER VALUE 
		P_SIGOUT			:	OUT	STD_LOGIC							-- FINAL SIGNAL BIT VALUE AFTER THE FILTER FUNCTION AND HYSTERISIS HAVE BEEN APPLIED

	);
END COMPONENT;

-- RS-485 SERIAL RECEIVE MODULE
COMPONENT SERIAL_RX is
port (
		MASTER_RST_B		:	IN	STD_LOGIC;							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
		CLK_5M_GL			:	IN	STD_LOGIC;
		RX_INPUT			:	IN	STD_LOGIC;							-- FINAL RX SIGNAL BIT STREAM AFTER THE FILTER FUNCTION AND HYSTERISIS HAVE BEEN APPLIED
		MODULE_ADDR			:	IN	STD_LOGIC_VECTOR(4 DOWNTO 0);		-- HARDWIRED ADDRESS OF THIS MODULE
		
		RX_WORD				:	OUT	STD_LOGIC_VECTOR(14 DOWNTO 0);		-- FINAL RECEIVED RX WORD
		RX_ODD_PARITY		:	OUT	STD_LOGIC;							-- ODD PARITY FOR THE RX_WORD
		RX_PARITY_ERR		:	OUT	STD_LOGIC;							-- LATCHED VESRION OF THE LAST RX PARITY ERROR
		RX_STRB				:	OUT	STD_LOGIC							-- SINGLE CLOCK PULSE STRB INDICATES THE RX_WORD WAS UPDATED
	);
END COMPONENT;

-- RS-485 SERIAL TRANSMIT MODULE
COMPONENT SERIAL_TX is
port (
		MASTER_RST_B		:	IN	STD_LOGIC;							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
		CLK_5M_GL			:	IN	STD_LOGIC;
		TX_WORD				:	IN	STD_LOGIC_VECTOR(14 DOWNTO 0);		-- PARALLEL WORD TO BE TRANSMITTED (NOTE--BIT 15 IS ODD PARITY CALCULATED AS SERIAL TX IS SENT)
		TX_STRB				:	IN	STD_LOGIC;							-- SINGLE CLOCK PULSE STRB INDICATES NEW TX_WORD READY FOR TX
		
		P_TX_EN				:	OUT	STD_LOGIC;							-- SERIAL TX DRIVER ENABLE
		SER_TX_BIT			:	OUT	STD_LOGIC							-- TX BIT STREAM
	);
END COMPONENT;

-- MAIN COMMUNICATION AND SEQUENCER MOPDULE
COMPONENT MAIN_SEQUENCER is
port (
		MASTER_RST_B		:	IN	STD_LOGIC;							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
		CLK_5M_GL			:	IN	STD_LOGIC;							-- MASTER 5 MHZ CLOCK
		
		SIGOUT_VOP_UVL		:	IN	STD_LOGIC;							-- UNDER-VOLTAGE LOCKOUT FAILSAFE ('1' = V_OP_RAIL FELL BELOW THE THRESHOLD)
				
		RECD_SER_WORD		:	IN	STD_LOGIC_VECTOR(14 DOWNTO 0);		-- WORD RECEIVED FROM THE SERIAL PORT
		SER_WORD_STB		:	IN	STD_LOGIC;							-- SINGLE CLOCK PULSE STROBE INDICATES AN UPDATED SERIAL WORD
		
		P_CH_MREG_EN_B		:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);		-- CHANNEL ENABLE SIGNAL: MAIN REGULATOR IC, ACTIVE LOW
		P_CH_IAUX_EN		:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);		-- CHANNEL ENABLE SIGNAL: IAUX REGULATOR IC, ACTIVE HIGH
		P_CH_VOSG_EN		:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);		-- CHANNEL ENABLE SIGNAL: VOS_GEN REGULATOR IC, ACTIVE HIGH
		
		P_COMPLETED_SEQ		:	OUT	STD_LOGIC;							-- PULSE INDICATES MAIN SEQUNEC COMPLETED
		
		CH_ACTIVE_STAT		:	OUT	STD_LOGIC							-- '1' INDICATES AT LEAST ONE CHANNEL ACTIVE
	);
END COMPONENT;

--===========SPECIAL TEST COMPONENTS:==============
COMPONENT SLOW_PULSE_EN_GEN is
port 	(
    		CLK_5M_GL		:	IN	STD_LOGIC;							-- FPGA MASTER CLOCK--ASSUMED TO BE 5 MHZ
    		MASTER_RST_B	:	IN	STD_LOGIC;							-- ACTIVE LOW RESET
			CNT_EN			:	IN	STD_LOGIC;							-- ACTIVE HIGH COUNT ENABLE
			SIM_10KX		:	IN	STD_LOGIC;							-- SPECIAL SIM MODE--SPEEDS UP BY 100,000 TIMES (1SEC=10USEC)

    		ONE_SEC_CLK_EN	:	OUT	STD_LOGIC							-- OUTPUT PULSE SIGNIFIES 1 SEC INTERVAL--SUITABLE FOR USE AS A CLOCK ENABLE.
		);
END COMPONENT;
		
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE INTERNAL SIGNALS
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

SIGNAL	MASTER_RST_B					:	STD_LOGIC;									-- POR_FPGA SYNC'D TO THE 40 MHZ CLOCK
SIGNAL	DEL0_DEV_RST_B					:	STD_LOGIC;									-- SYNC FF FOR FOR GENERATING THE MASTER_RST_B

SIGNAL	CLK_5M_GL, N_CLK_5M_GL			:	STD_LOGIC;									-- GENERATED 5 MHZ CLOCK--MASTER CLOCK!!!!
SIGNAL	REFCNT, N_REFCNT				:	INTEGER RANGE 0 TO 3;						-- COUNTER USED TO GENERATE THE CLK_5M_GL

SIGNAL	RS485_RX1_IN, RS485_RX0_IN		:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- USED TO SYNC RX_SIG_IN TO THE 5MHZ CLOCK
SIGNAL	FILTD_RS485RX					:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- FILTERED RX SIGNAL FOR THE RS-485 PORT

SIGNAL	UVL_VOP0_IN, UVL_VOP_FILT_IN	:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- USED TO SYNC UVL_VOP_IN TO THE 5MHZ CLOCK
SIGNAL	LAT_VOP_UVL, N_LAT_VOP_UVL		:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- LATCHED COPY OF THE VOP UVL---CLEARED BY THE 1 HZ TX STRB

SIGNAL  ENABLES_SEU_DET, N_ENABLES_SEU_DET	:	STD_LOGIC_VECTOR(0 DOWNTO 0);			-- LATCHED VESRION OF THE SEU DETECT FOR THE 24 ENABLES.

SIGNAL	UVL_1V5_0IN, UVL_1V5_1IN		:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- USED TO SYNC UVL_1V5_IN TO THE 5MHZ CLOCK
SIGNAL	LAT_1V5_UVL, N_LAT_1V5_UVL		:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- LATCHED COPY OF THE 1V5 UVL---CLEARED BY THE 1 HZ TX STRB

SIGNAL 	CH_EN_0SIG, CH_EN_1SIG			:	STD_LOGIC_VECTOR(7 DOWNTO 0);				-- USED TO SYNC EXT_CH_EN_PORT TO THE 5 MHZ CLOCK

SIGNAL	FILTD_TEMP_OK_B					:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- FILTERED VERSION OF TEMP_OK_B
SIGNAL	FILTD_FUSE_1_2_OK				:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- FILTERED VERSION OF FUSE_1_2_OK UVL INPUT
SIGNAL	FILTD_FUSE_3_4_OK				:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- FILTERED VERSION OF FUSE_3_4_OK UVL INPUT
SIGNAL	FILTD_FUSE_5_6_OK				:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- FILTERED VERSION OF FUSE_5_6_OK UVL INPUT
SIGNAL	FILTD_FUSE_7_8_OK				:	STD_LOGIC_VECTOR(0 DOWNTO 0);				-- FILTERED VERSION OF FUSE_7_8_OK UVL INPUT

SIGNAL	FILT_SIGOUT_RX					: 	STD_LOGIC_VECTOR(7 DOWNTO 0);				-- FINAL OUTPUT SIGNAL FILTER VALUE FOR THE RX RECEIVE (FOR SIM DEBUG)
SIGNAL	SIGOUT_RX						:	STD_LOGIC;									-- FINAL SIGNAL OUT AFTER FILTER AND HYSTERISIS APPLIED

SIGNAL	FILT_VOPOUT_UVL					: 	STD_LOGIC_VECTOR(7 DOWNTO 0);				-- FINAL OUTPUT SIGNAL FILTER VALUE FOR THE VOP UVL (FOR SIM DEBUG)
SIGNAL	SIGOUT_VOP_UVL					:	STD_LOGIC;									-- FINAL SIGNAL OUT AFTER FILTER AND HYSTERISIS APPLIED

SIGNAL	RX_WORD							:	STD_LOGIC_VECTOR(14 DOWNTO 0);				-- RECEIVED SERIAL WORD BUFFER
SIGNAL	RX_STRB							:	STD_LOGIC;									-- STROBE PULSE, 1 CLOCK WIDE, INDICATES NEW RX WORD READY
SIGNAL	RX_ODD_PARITY					:	STD_LOGIC;									-- ODD PARITY BIT FOR RX WORD (FOR SIM DEBUG)
SIGNAL	RX_PARITY_ERR					:	STD_LOGIC;									-- LATCHED VERSION OF THE LAST RX ODD PARITY ERROR

SIGNAL	TEST_TX_STROBE					:	STD_LOGIC;	
SIGNAL	SERIAL_TX_BIT					:	STD_LOGIC;
SIGNAL	SER_TX_EN						:	STD_LOGIC;									-- SERIAL TX DRIVER ENABLE

CONSTANT	UPPER_HYS_THRESH			:	STD_LOGIC_VECTOR(7 DOWNTO 0) := "01001100";	-- UPPER HYSTERISIS THRESHOLD = 76 COUNTS OF 255 (ACTUALLY 240 WITH TRUNCATION EFFECTS)
CONSTANT	LOWER_HYS_THRESH			:	STD_LOGIC_VECTOR(7 DOWNTO 0) := "00101100";	-- UPPER HYSTERISIS THRESHOLD =  44 COUNTS OF 255 (ACTUALLY 240 WITH TRUNCATION EFFECTS)

SIGNAL 	CH_MREG_EN_B					:	STD_LOGIC_VECTOR(7 DOWNTO 0);				-- CHANNEL ENABLE SIGNAL: MAIN REGULATOR IC, ACTIVE LOW
SIGNAL	CH_IAUX_EN						:	STD_LOGIC_VECTOR(7 DOWNTO 0);				-- CHANNEL ENABLE SIGNAL: IAUX REGULATOR IC, ACTIVE HIGH
SIGNAL	CH_VOSG_EN						:	STD_LOGIC_VECTOR(7 DOWNTO 0);				-- CHANNEL ENABLE SIGNAL: VOS_GEN REGULATOR IC, ACTIVE HIGH

-- FOR SPECIAL TEST MUX SUPPORT--NEED REGISTER TO AVOID GLITCHES
SIGNAL 	N_MUX_CH_MREG_EN_B, MUX_CH_MREG_EN_B	:	STD_LOGIC_VECTOR(7 DOWNTO 0);				-- CHANNEL ENABLE SIGNAL: MAIN REGULATOR IC, ACTIVE LOW
SIGNAL	N_MUX_CH_IAUX_EN, MUX_CH_IAUX_EN		:	STD_LOGIC_VECTOR(7 DOWNTO 0);				-- CHANNEL ENABLE SIGNAL: IAUX REGULATOR IC, ACTIVE HIGH
SIGNAL	N_MUX_CH_VOSG_EN, MUX_CH_VOSG_EN		:	STD_LOGIC_VECTOR(7 DOWNTO 0);				-- CHANNEL ENABLE SIGNAL: VOS_GEN REGULATOR IC, ACTIVE HIGH

SIGNAL 	CH_ACTIVE_STAT					:	STD_LOGIC;									-- '1' INDICATES AT LEAST ONE CHANNEL ACTIVE

SIGNAL TRANSMIT_WORD, N_TRANSMIT_WORD	:	STD_LOGIC_VECTOR(15 DOWNTO 0);				-- PARALLEL WORD TO BE TRANSMITTED (NOTE--BIT 15 IS ODD PARITY CALCULATED AS SERIAL TX IS SENT)

SIGNAL COMPLETED_MAIN_SEQ				:	STD_LOGIC;									-- PULSE INDICATES THAT THE MAIN SEQUENCE COMPLETED

SIGNAL	N_PREV_RX_WORD, PREV_RX_WORD	:	STD_LOGIC_VECTOR(14 DOWNTO 0); 				-- LATCHED COPY OF THE LAST SERIAL RX WORD MODULO 2 BITS

SIGNAL	N_PREV_EN_STATE, PREV_EN_STATE	:	STD_LOGIC_VECTOR(23 DOWNTO 0);				-- SAVED COPY OF THE 24 ENABLE BITS USED FOR COMPARISON

SIGNAL	N_PREV_RX_PARITY_ERR, PREV_RX_PARITY_ERR	:	STD_LOGIC;						-- SAVED COPY OF THE RX PARITY ERROR

-- DIP SWITCH OVERRIDE REGISTER:  THIS REGISTER CAN ONLY WRITE TO ONE BIT AT A TIME.  BOTH BITS MUST BE '1' TO BE IN OVERRIDE MODE.  THEREFORE 2 SUCCESSIVE WRITES ARE NEEDED.
-- EXAMPLE:  '01' FOLLOWED BY '11' 
SIGNAL	SW_OVERRIDE						:	STD_LOGIC_VECTOR(1 DOWNTO 0);				-- '11' = OVERRIDE MODE.  ALL OTHER STATES = NORMAL SWITCH MODE DRIVEN OPERATION


--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- TEMPORARY PLACEHOLDERS!!!!!!!!!

SIGNAL MAN_GPIO_ENABLES					:	STD_LOGIC_VECTOR(0 DOWNTO 0):= "0";			-- ENABLES MANUAL GPIO PORT---AKA MASTER_SLAVEB_SEL FOR SPECIAL THIS TEST VERSION



--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
BEGIN
-- THIS PROCESS SYNCHRONIZES THE EXTERNAL POR_FPGA SIGNAL TO THE 40 MHZ CLOCK
SYNC_DEV_RST_B:PROCESS(POR_FPGA, CLK40M_OSC)
    BEGIN
        IF POR_FPGA = '0' THEN
			DEL0_DEV_RST_B		<=	'0';
			MASTER_RST_B		<=	'0';
		
        ELSIF (CLK40M_OSC'EVENT AND CLK40M_OSC='1') THEN
			DEL0_DEV_RST_B		<=	POR_FPGA;
			MASTER_RST_B		<=	DEL0_DEV_RST_B;
		
        END IF;

    END PROCESS SYNC_DEV_RST_B;
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- REGISTERS USED TO GENERATE A 5 MHZ CLOCK (DIV-BY-4 FOLLOWED BY DIV-BY-2)
GENCLKREG:PROCESS(MASTER_RST_B, CLK40M_OSC)
    BEGIN
        IF MASTER_RST_B = '0' THEN
			CLK_5M_GL	<=	'0';
			REFCNT		<=	 0;
		
        ELSIF (CLK40M_OSC'EVENT AND CLK40M_OSC='1') THEN
			CLK_5M_GL	<=	N_CLK_5M_GL;
			REFCNT		<=	N_REFCNT;

        END IF;

    END PROCESS GENCLKREG;

-- PROCESS TO GENERATE THE 5 MHZ CLOCK
GEN_5M_CLK:PROCESS(REFCNT, CLK_5M_GL)
	BEGIN
		IF REFCNT > 2 THEN
			N_REFCNT		<=	0;
			N_CLK_5M_GL		<=	NOT(CLK_5M_GL);
			
		ELSE
			N_REFCNT		<=	REFCNT + 1;
			N_CLK_5M_GL		<=	CLK_5M_GL;
		END IF;
	END PROCESS;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE ALL REGISTERS THAT USE THE 5 MHZ CLOCK
REG5M:PROCESS(CLK_5M_GL, MASTER_RST_B)	
	BEGIN
		IF MASTER_RST_B = '0' THEN
			RS485_RX0_IN	<=	 "0";										-- CLK SYNCHRONIZING REGISTER
			RS485_RX1_IN	<=	 "0";										-- CLK SYNCHRONIZING REGSITER

			UVL_VOP0_IN		<=	 "0";										-- CLK SYNCHRONIZING REGISTER
			UVL_VOP_FILT_IN	<=	 "0";										-- CLK SYNCHRONIZING REGSITER 
			LAT_VOP_UVL		<=	 "0";										-- LATCHED VERSION

			UVL_1V5_0IN		<=	 "0";										-- CLK SYNCHRONIZING REGISTER
			UVL_1V5_1IN		<=	 "0";										-- CLK SYNCHRONIZING REGISTER
			LAT_1V5_UVL		<=	 "0";										-- LATCHED VERSION

			
			CH_EN_0SIG		<=	 (OTHERS => '0');							-- CLK SYNCHRONIZING REGSITER
			CH_EN_1SIG		<=	 (OTHERS => '0');							-- CLK SYNCHRONIZING REGSITER
			
			TRANSMIT_WORD	<=	(OTHERS => '0');
			
			MUX_CH_MREG_EN_B	<=	(OTHERS => '0');						-- SPECIAL TEST SUPPORT REGISTERED MUX
			MUX_CH_IAUX_EN		<=	(OTHERS => '0');						-- SPECIAL TEST SUPPORT REGISTERED MUX
			MUX_CH_VOSG_EN		<=	(OTHERS => '0');						-- SPECIAL TEST SUPPORT REGISTERED MUX
			
			ENABLES_SEU_DET	<=	(OTHERS => '0');	
			PREV_EN_STATE	<=	(OTHERS => '0');
			
			PREV_RX_PARITY_ERR	<=	'0';
			
			PREV_RX_WORD		<=	(OTHERS => '0');

			
		ELSIF (CLK_5M_GL'EVENT AND CLK_5M_GL='1') THEN
			RS485_RX0_IN	<=	RX_FPGA;
			RS485_RX1_IN	<=	RS485_RX0_IN;								-- INPUT SIGNAL FULLY SYNC'D TO 5 MHZ CLOCK

			UVL_VOP0_IN		<=	UVL_VOP_IN;
			UVL_VOP_FILT_IN	<=	UVL_VOP0_IN;								-- INPUT SIGNAL FULLY SYNC'D TO 5 MHZ CLOCK
			LAT_VOP_UVL		<=	N_LAT_VOP_UVL;								-- LATCHED VERSION OF THE FILTERED VOP UVL SIGNAL

			UVL_1V5_0IN		<=	UVL_1V5_IN;
			UVL_1V5_1IN		<=	UVL_1V5_0IN;
			LAT_1V5_UVL		<=	N_LAT_1V5_UVL;								-- LATCHED VERSION OF THE UNFILTERED, BUT SYNC'D VERSION OF THE 1V5 UVL
			
			CH_EN_0SIG		<=	EXT_CH_EN_PORT;
			CH_EN_1SIG		<=	CH_EN_0SIG;									-- INPUT SIGNAL FULLY SYNC'D TO 5 MHZ CLOCK
			
			TRANSMIT_WORD	<=	N_TRANSMIT_WORD;

			MUX_CH_MREG_EN_B	<=	N_MUX_CH_MREG_EN_B;						-- SPECIAL TEST SUPPORT REGISTERED MUX
			MUX_CH_IAUX_EN		<=	N_MUX_CH_IAUX_EN;						-- SPECIAL TEST SUPPORT REGISTERED MUX
			MUX_CH_VOSG_EN		<=	N_MUX_CH_VOSG_EN;						-- SPECIAL TEST SUPPORT REGISTERED MUX
			
			ENABLES_SEU_DET	<=	N_ENABLES_SEU_DET;
			PREV_EN_STATE	<=	N_PREV_EN_STATE;
			
			PREV_RX_PARITY_ERR	<=	N_PREV_RX_PARITY_ERR;
			
			PREV_RX_WORD	<=	N_PREV_RX_WORD;
		END IF;
		
	END PROCESS;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- placeholder
-- PROCESS THAT WAITS FOR >35 '0' BITS FOLLOWED BY 2 START BITS IN THE FILTERED RS485 RX LINE AND THEN GENERATES 36 CLOCK CYCLES 



--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- placeholder
-- PROCESS THAT PERFORMS THE MUX SELECTION OF EITHER THE RS485 OR THE SPI POR CLOCK AND SERIAL DATA SOURCES 



--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

-- APPEARS THAT A LOT OF REWORK IS NEEDED FOR THIS PROCESS TO REMOVE THE OLD SPECIAL TEST FEATURES!!!!

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- PROCESS THE STATUS BITS FOR BOTH TX AND RX :
-- (1) MUXES THE 4 BIT STATUS OUTPUT SENT TO MUX FPGA PINS WHEN USED AS A MASTER OUTPUT FUNCTION (VERSUS NORMAL SLAVE OUTPUT ENABLES)
-- (2) CONCATINATES AND LATCHES A COPY OF WORD TO BE TRANSMITTED (USED BY SLAVE TO COLLECT STATUS OF IRRADIATED BOARD)
-- (3) LATCHES DETECTED CHANGES IN THE UVL BITS DURING THE ENTIRE PERIOD BETWEEN TRANSMIT PULSE TRIGGERS
-- (4) LATCHES DETECTED CHANGES IN THE 24 ENABLE BITS DURING THE ENTIRE PERIOD BETWEEN TRANSMIT PULSE TRIGGERS

-- NOTE:	SIGOUT_VOP_UVL USES IIR FILTER, BUT UVL_1V5_1IN DOES NOT.  THIS IS BECAUSE THE FPGA IS NOT OPERATING IF UVL_1V5_1IN IS ACTIVE
-- 			SINCE THIS IS NORMALLY A HARDWIRED FAILSAFE.  IT IS BEING BROUGHT OUT HERE FOR THIS SPECIAL TEST CONFIG.
-- CH_EN_1SIG:  	X8 EXTERNAL GPIO JUMPERS 
-- UVL_BITS: 		X2 BITS FOR THE 1V5 AND VOP UVL SIGNALS
-- ADDR_SEL:		X5 MODULE ADDRESS JUMPER BITS 
-- SIGOUT_VOP_UVL:	X1 UVL FOR THE VOP RAIL (FILTERED USING THE IIR MODULE)
-- UVL_1V5_1IN:		X1 UVL FOR THE 1V5 RAIL (ONLY SYNC'S TO THE 5 MHZ CLOCK---NOT FILTERED)
--		RX_WORD:	EN_SEU & UVL_BITS & ADDR_SEL & CH_EN_1SIG;

-- NOTE: MAN_GPIO_ENABLES == MASTER_SLAVEB_SEL FOR THIS SPECIAL TEST VERSION

STATUS:PROCESS(		RX_WORD, RX_STRB, MAN_GPIO_ENABLES, RX_PARITY_ERR, UVL_1V5_1IN, SIGOUT_VOP_UVL, ENABLES_SEU_DET, TRANSMIT_WORD, LAT_VOP_UVL, LAT_1V5_UVL,
					CH_VOSG_EN, CH_IAUX_EN, CH_MREG_EN_B, TEST_TX_STROBE, PREV_RX_PARITY_ERR,
					CH_EN_1SIG, PREV_RX_WORD, ADDR_SEL, PREV_EN_STATE
				)
	BEGIN
	
-- ++++++++  LATCH UVL SIGNALS HERE  ++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
		IF 		UVL_1V5_1IN = "1" 		THEN									-- LATCH ANY DETECTED CHANGE IN THE 1V5 UVL BIT STATE
					N_LAT_1V5_UVL	<=	"1";
		ELSIF 	TEST_TX_STROBE = '1'	THEN									-- LATCHED STATE CLEARED ONCE READ BY THE TX MODULE (SEE BELOW)
					N_LAT_1V5_UVL 	<=	"0";
		ELSE
					N_LAT_1V5_UVL 	<=  LAT_1V5_UVL;
		END IF;
		
		
		IF 		SIGOUT_VOP_UVL = '1' 	THEN									-- LATCH ANY DETECTED CHANGE IN THE VOP UVL BIT STATE
					N_LAT_VOP_UVL	<=	"1";
		ELSIF 	TEST_TX_STROBE = '1'	THEN									-- LATCHED STATE CLEARED ONCE READ BY THE TX MODULE (SEE BELOW)
					N_LAT_VOP_UVL 	<=	"0";
		ELSE
					N_LAT_VOP_UVL 	<=	LAT_VOP_UVL;
		END IF;	

-- ++++++++  LATCH SEU DETECTION BIT OF 24 ENABLE SIGNALS HERE  +++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
		IF TEST_TX_STROBE = '1' 		THEN
			N_PREV_EN_STATE	<=	CH_MREG_EN_B & CH_IAUX_EN & CH_VOSG_EN;			-- SAVE A COPY OF ALL 24 ENABLE BITS
		ELSE
			N_PREV_EN_STATE	<=	PREV_EN_STATE;
		END IF;
	
		IF 		PREV_EN_STATE	/= CH_MREG_EN_B & CH_IAUX_EN & CH_VOSG_EN THEN	-- SET THE BIT IS THE NOT EQUAL CONDITION DETECTED
					N_ENABLES_SEU_DET		<=	"1";
		ELSIF 	TEST_TX_STROBE = '1' 	THEN									-- ONLY CLEAR THE BIT ONCE READ FOR TX
					N_ENABLES_SEU_DET		<=	"0";
		ELSE
					N_ENABLES_SEU_DET		<=	ENABLES_SEU_DET;
		END IF;
		
-- ++++++++  CONCATINATE AND STORE A COPY OF THE TX WORD HERE	(SEE DESCRIPTIONS ABOVE)+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
		IF TEST_TX_STROBE = '1'	THEN
			N_TRANSMIT_WORD		<=	ENABLES_SEU_DET & LAT_VOP_UVL & LAT_1V5_UVL & ADDR_SEL(4 DOWNTO 0) & CH_EN_1SIG(7 DOWNTO 0);
		ELSE
			N_TRANSMIT_WORD		<=	TRANSMIT_WORD;
		END IF;

-- ++++++++  MUX SIGNALS OF RX DATA HERE  ++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++		
		IF RX_STRB = '1' 		THEN
			N_PREV_RX_WORD					<=	RX_WORD;
			N_PREV_RX_PARITY_ERR			<=	RX_PARITY_ERR;
		ELSE
			N_PREV_RX_WORD					<=	PREV_RX_WORD;
			N_PREV_RX_PARITY_ERR			<=	PREV_RX_PARITY_ERR;
		END IF;

		IF MAN_GPIO_ENABLES = "1"	THEN	
			N_MUX_CH_MREG_EN_B(0)			<=	PREV_RX_PARITY_ERR;							-- DETECTED PARITY ERROR STATE
			N_MUX_CH_IAUX_EN(0)				<=	PREV_RX_WORD(14);							-- ENABLE SEU FLIP DETECTED
			N_MUX_CH_VOSG_EN(0)				<=	PREV_RX_WORD(12);							-- 1V5 UVL STATUS

			N_MUX_CH_MREG_EN_B(1)			<=	PREV_RX_WORD(13);							-- VOP UVL STATUS
			N_MUX_CH_IAUX_EN(1)				<=	'0';
			N_MUX_CH_VOSG_EN(1)				<=	'0';
		
			N_MUX_CH_MREG_EN_B(7 DOWNTO 2)	<=	(OTHERS => '0');
			N_MUX_CH_IAUX_EN(7 DOWNTO 2)	<=	(OTHERS => '0');
			N_MUX_CH_VOSG_EN(7 DOWNTO 2)	<=	(OTHERS => '0');
			
		ELSE
			N_MUX_CH_MREG_EN_B(7 DOWNTO 0)	<=	CH_MREG_EN_B(7 DOWNTO 0);
			N_MUX_CH_IAUX_EN(7 DOWNTO 0)	<=	CH_IAUX_EN(7 DOWNTO 0);
			N_MUX_CH_VOSG_EN(7 DOWNTO 0)	<=	CH_VOSG_EN(7 DOWNTO 0);
			
		END IF;

	END PROCESS;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- INSTANTIATE THE IIR FILTER COMPONENT FOR THE SERIAL RECEIVE SIGNAL OF THE RS485 INTERFACE
RS485_RX_FILT:IIR_FILT
port MAP(
			MASTER_RST_B		=>	MASTER_RST_B,							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
			CLK_5M_GL			=>	CLK_5M_GL,								-- MASTER 5 MHZ CLOCK
			
			SIG_IN				=>	RS485_RX1_IN,							-- RS-485 SIGNAL TO BE FILTERED
			THRESH_UPPER		=>	UPPER_HYS_THRESH,						-- UPPER HYSTERISIS THRESHOLD (IE RISING SIGNAL THRESHOLD)
			THRESH_LOWER		=> 	LOWER_HYS_THRESH,						-- LOWER HYSTERISIS THRESHOLD (IE FALLING SIGNAL THRESHOLD)
			FILT_SIGOUT			=>	FILT_SIGOUT_RX,							-- SIGNAL FILTER OUTPUT VALUE FOR THE RX SIGNAL
			P_SIGOUT			=>	FILTD_RS485RX							-- FINAL SIGNAL BIT VALUE AFTER THE FILTER FUNCTION AND HYSTERISIS HAVE BEEN APPLIED

		);
		
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- INSTANTIATE THE IIR FILTER COMPONENT FOR THE VOP UNDERVOLTAGE LOCKOUT SIGNAL
VOP_UVL_FILT:IIR_FILT
port MAP(
			MASTER_RST_B		=>	MASTER_RST_B,							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
			CLK_5M_GL			=>	CLK_5M_GL,								-- MASTER 5 MHZ CLOCK
			
			SIG_IN				=>	UVL_VOP_FILT_IN,						-- SIGNAL TO BE FILTERED
			THRESH_UPPER		=>	UPPER_HYS_THRESH,						-- UPPER HYSTERISIS THRESHOLD (IE RISING SIGNAL THRESHOLD)
			THRESH_LOWER		=> 	LOWER_HYS_THRESH,						-- LOWER HYSTERISIS THRESHOLD (IE FALLING SIGNAL THRESHOLD)
			FILT_SIGOUT			=>	FILT_VOPOUT_UVL,						-- SIGNAL FILTER OUTPUT VALUE FOR THE RX SIGNAL
			P_SIGOUT			=>	SIGOUT_VOP_UVL							-- FINAL SIGNAL BIT VALUE AFTER THE FILTER FUNCTION AND HYSTERISIS HAVE BEEN APPLIED

		);

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- INSTANTIATE THE SERIAL RX MODULE		
SERIAL_REC:SERIAL_RX
port MAP (
			MASTER_RST_B		=>	MASTER_RST_B,							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
			CLK_5M_GL			=>	CLK_5M_GL,
			RX_INPUT			=>	SIGOUT_RX,									-- FINAL RX SIGNAL BIT STREAM AFTER THE FILTER FUNCTION AND HYSTERISIS HAVE BEEN APPLIED
			MODULE_ADDR			=>	ADDR_SEL,								-- ADDRESS FOR THIS MODULE
			
			RX_WORD				=>	RX_WORD,								-- FINAL RECEIVED RX WORD
			RX_ODD_PARITY		=>	RX_ODD_PARITY,							-- ODD PARITY FOR THE RX_WORD
			RX_PARITY_ERR		=>	RX_PARITY_ERR,							-- LATCHED VERSION OF THE LAST RX PARITY ERROR
			RX_STRB				=>	RX_STRB									-- SINGLE CLOCK PULSE STRB INDICATES THE RX_WORD WAS UPDATED
		);

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- INSTANTIATE THE SERIAL TX MODULE	COMPONENT
SERIAL_TRANS:SERIAL_TX
port MAP(
			MASTER_RST_B		=>	MASTER_RST_B,							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
			CLK_5M_GL			=>	CLK_5M_GL,
			TX_WORD				=>	TRANSMIT_WORD,							-- PARALLEL WORD TO BE TRANSMITTED (NOTE--BIT IS ODD PARITY CALCULATED AS SERIAL TX IS SENT)
			TX_STRB				=>	TEST_TX_STROBE,							-- SINGLE CLOCK PULSE STRB INDICATES NEW TX_WORD READY FOR TX
			
			P_TX_EN				=>	SER_TX_EN,								-- SERIAL TX DRIVER ENABLE
			SER_TX_BIT			=>	SERIAL_TX_BIT							-- TX BIT STREAM
	);

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- INSTANTIATE THE MAIN COMMUNICATIONS AND SEQUENCER MODULE
CONTROL:MAIN_SEQUENCER
port MAP (
			MASTER_RST_B		=>	MASTER_RST_B,							-- RESET WITH ASYNC ASSERT, BUT SYNCHRONIZED TO THE 40 MHZ CLOCK EDGE
			CLK_5M_GL			=>	CLK_5M_GL,								-- MASTER 5 MHZ CLOCK
			
			SIGOUT_VOP_UVL		=>	SIGOUT_VOP_UVL,							-- UNDER-VOLTAGE LOCKOUT ('1' = V_OP_RAIL FELL BELOW THE THRESHOLD)
					
			RECD_SER_WORD		=>	RX_WORD,								-- WORD RECEIVED FROM THE SERIAL PORT
			SER_WORD_STB		=>	RX_STRB,								-- SINGLE CLOCK PULSE STROBE INDICATES AN UPDATED SERIAL WORD
			
			P_CH_MREG_EN_B		=>	CH_MREG_EN_B,							-- CHANNEL ENABLE SIGNAL: MAIN REGULATOR IC, ACTIVE LOW
			P_CH_IAUX_EN		=>	CH_IAUX_EN,								-- CHANNEL ENABLE SIGNAL: IAUX REGULATOR IC, ACTIVE HIGH
			P_CH_VOSG_EN		=>	CH_VOSG_EN,								-- CHANNEL ENABLE SIGNAL: VOS_GEN REGULATOR IC, ACTIVE HIGH
			
			P_COMPLETED_SEQ		=>	COMPLETED_MAIN_SEQ,						-- PULSE INDICATES SEQUENCE COMPLETED
			
			CH_ACTIVE_STAT		=> 	CH_ACTIVE_STAT							-- '1' INDICATES AT LEAST ONE CHANNEL ACTIVE
		);

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- INSTANTIATE A 1 HZ PULSE GENERATOR USED FOR SPECIAL TEST TO STRB THE TX FUNCTION 		
TX_PROMPT:SLOW_PULSE_EN_GEN
port MAP (
    		CLK_5M_GL			=>	CLK_5M_GL,								-- FPGA MASTER CLOCK--ASSUMED TO BE 5 MHZ
    		MASTER_RST_B		=>	MASTER_RST_B,							-- ACTIVE LOW RESET
			CNT_EN				=>	'1',									-- ACTIVE HIGH COUNT ENABLE
			SIM_10KX			=>	'0',									-- SPECIAL SIM MODE--SPEEDS UP  (1SEC=1000USEC)

    		ONE_SEC_CLK_EN		=>	TEST_TX_STROBE							-- OUTPUT PULSE SIGNIFIES 1 SEC INTERVAL--SUITABLE FOR USE AS A CLOCK ENABLE.
		);
		
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- ASSIGN INTERNAL SIGNALS TOP EXTERNAL PORTS
P_MASTER_RST_B		<=	MASTER_RST_B;
P_CLK_5M_GL			<=	CLK_5M_GL;

P_CH_MREG_EN_B		<=	MUX_CH_MREG_EN_B;							-- CHANNEL ENABLE SIGNAL: MAIN REGULATOR IC, ACTIVE LOW
P_CH_IAUX_EN		<=	MUX_CH_IAUX_EN;								-- CHANNEL ENABLE SIGNAL: IAUX REGULATOR IC, ACTIVE HIGH
P_CH_VOSG_EN		<=	MUX_CH_VOSG_EN;								-- CHANNEL ENABLE SIGNAL: VOS_GEN REGULATOR IC, ACTIVE HIGH
CH_STAT_LED			<=	CH_ACTIVE_STAT;

P_SERIAL_TX			<=	CONV_STD_LOGIC_VECTOR(SERIAL_TX_BIT, 1);

P_SER_TX_EN			<=	'1';										-- LEAVING STUCK ON FOR TEST,,,,WAS SER_TX_EN;

TX_EN				<=	"0";										-- LEAVING STUCK OFF AS RX FOR TEST 

end RTL;